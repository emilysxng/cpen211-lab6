//cpu testbench here